//Verilog HDL for "MultiChannel_EMG_Model", "MultiChannelAFE_TB" "functional"


module MultiChannelAFE_TB ( );

endmodule
